class apb_test_rd_cmd_seq;
    apb_env env;
    virtual apb_if vif;

    
endclass
